library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

use work.Types.all;

package SramPack is
  constant SramDataW : positive := 16;
  constant SramAddrW : positive := 18;

end package;

package body SramPack is

end package body;
 
